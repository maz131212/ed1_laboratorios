///// ELECTRÓNICA DIGITAL 1
///// AXEL MAZARIEGOS - 131212
///// 31 - OCTUBRE - 2020
/////
///// LABORATORIO 09
///// EJERCICIO 05



module  ROM(input wire  [6:0] A,
            output reg  [12:0] Y);


  always @(A)
  begin

    if (A[0])

      casez (A) //casez para que reconozca los don't care
        7'b00001?1 : Y <= 13'b0100000001000;
        7'b00000?1 : Y <= 13'b1000000001000;
        7'b00011?1 : Y <= 13'b1000000001000;
        7'b00010?1 : Y <= 13'b0100000001000;
        7'b0010??1 : Y <= 13'b0001001000010;
        7'b0011??1 : Y <= 13'b1001001100000;
        7'b0100??1 : Y <= 13'b0011010000010;
        7'b0101??1 : Y <= 13'b0011010000100;
        7'b0110??1 : Y <= 13'b1011010100000;
        7'b0111??1 : Y <= 13'b1000000111000;
        7'b1000?11 : Y <= 13'b0100000001000;
        7'b1000?01 : Y <= 13'b1000000001000;
        7'b1001?11 : Y <= 13'b1000000001000;
        7'b1001?01 : Y <= 13'b0100000001000;
        7'b1010??1 : Y <= 13'b0011011000010;
        7'b1011??1 : Y <= 13'b1011011100000;
        7'b1100??1 : Y <= 13'b0100000001000;
        7'b1101??1 : Y <= 13'b0000000001001;
        7'b1110??1 : Y <= 13'b0011100000010;
        7'b1111??1 : Y <= 13'b1011100100000;
        default : Y =13'b0000000000000;

        endcase

      else Y <= 13'b1000000001000;

  end

endmodule





// este fue un modulo hecho escribiendo todoas las posibles combinaciones
// sin utilizar don't cares
/*module  ROM(input wire  [6:0] A,
            output reg  [12:0] Y);


  always @(A)
  begin

    if (A[0])

      case (A)
        7'b0000101 : Y <= 13'b0100000001000;
        7'b0000111 : Y <= 13'b0100000001000;

        7'b0000001 : Y <= 13'b1000000001000;
        7'b0000011 : Y <= 13'b1000000001000;

        7'b0001101 : Y <= 13'b1000000001000;
        7'b0001111 : Y <= 13'b1000000001000;

        7'b0001001 : Y <= 13'b0100000001000;
        7'b0001011 : Y <= 13'b0100000001000;

        7'b0010001 : Y <= 13'b0001001000010;
        7'b0010011 : Y <= 13'b0001001000010;
        7'b0010101 : Y <= 13'b0001001000010;
        7'b0010111 : Y <= 13'b0001001000010;

        7'b0011001 : Y <= 13'b1001001100000;
        7'b0011011 : Y <= 13'b1001001100000;
        7'b0011101 : Y <= 13'b1001001100000;
        7'b0011111 : Y <= 13'b1001001100000;

        7'b0100001 : Y <= 13'b0011010000010;
        7'b0100011 : Y <= 13'b0011010000010;
        7'b0100101 : Y <= 13'b0011010000010;
        7'b0100111 : Y <= 13'b0011010000010;

        7'b0101001 : Y <= 13'b0011010000100;
        7'b0101011 : Y <= 13'b0011010000100;
        7'b0101101 : Y <= 13'b0011010000100;
        7'b0101111 : Y <= 13'b0011010000100;

        7'b0110001 : Y <= 13'b1011010100000;
        7'b0110011 : Y <= 13'b1011010100000;
        7'b0110101 : Y <= 13'b1011010100000;
        7'b0110111 : Y <= 13'b1011010100000;

        7'b0111001 : Y <= 13'b1000000111000;
        7'b0111011 : Y <= 13'b1000000111000;
        7'b0111101 : Y <= 13'b1000000111000;
        7'b0111111 : Y <= 13'b1000000111000;

        7'b1000011 : Y <= 13'b0100000001000;
        7'b1000111 : Y <= 13'b0100000001000;

        7'b1000001 : Y <= 13'b1000000001000;
        7'b1000101 : Y <= 13'b1000000001000;

        7'b1001011 : Y <= 13'b1000000001000;
        7'b1001111 : Y <= 13'b1000000001000;

        7'b1001001 : Y <= 13'b0100000001000;
        7'b1001101 : Y <= 13'b0100000001000;

        7'b1010001 : Y <= 13'b0011011000010;
        7'b1010011 : Y <= 13'b0011011000010;
        7'b1010101 : Y <= 13'b0011011000010;
        7'b1010111 : Y <= 13'b0011011000010;

        7'b1011001 : Y <= 13'b1011011100000;
        7'b1011011 : Y <= 13'b1011011100000;
        7'b1011101 : Y <= 13'b1011011100000;
        7'b1011111 : Y <= 13'b1011011100000;
        
        7'b1100001 : Y <= 13'b0100000001000;
        7'b1100011 : Y <= 13'b0100000001000;
        7'b1100101 : Y <= 13'b0100000001000;
        7'b1100111 : Y <= 13'b0100000001000;
        
        7'b1101001 : Y <= 13'b0000000001001;
        7'b1101011 : Y <= 13'b0000000001001;
        7'b1101101 : Y <= 13'b0000000001001;
        7'b1101111 : Y <= 13'b0000000001001;
        
        7'b1110001 : Y <= 13'b0011100000010;
        7'b1110011 : Y <= 13'b0011100000010;
        7'b1110101 : Y <= 13'b0011100000010;
        7'b1110111 : Y <= 13'b0011100000010;

        7'b1111001 : Y <= 13'b1011100100000;
        7'b1111011 : Y <= 13'b1011100100000;
        7'b1111101 : Y <= 13'b1011100100000;
        7'b1111111 : Y <= 13'b1011100100000;

        default : Y =13'b0000000000000;

        endcase

      //cuando el bit menos signifcativo es 0
      else Y <= 13'b1000000001000; 

  end

endmodule */


